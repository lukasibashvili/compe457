module mux_y(
  input [31:0] Ard,
  input [3:0] jump,
  input select,
  output [31:0] out
);

  always @(*)begin

    //keep it simple, how did you come up with smth like that?

  end

endmodule
