module mux_src1(
  input [31:0] Rn,
  input [31:0] Rs,
  input [31:0] PC_out,
  input [1:0] select,
  output [31:0] out
);

  always @(*)begin

    //rewrite as case statement

  end

endmodule
